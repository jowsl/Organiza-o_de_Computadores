module questao3 (s, maquina, out);
    input[2:0]s;


endmodule